module cla4(a, b, ci, co, s);
	input [3:0] a, b;
	input ci;
	output co;
	output [3:0] s;
	wire [2:0] c;
	
	// connect with 4 full adders which have no carry out
	fa_v2 cla_fa0 (.a(a[0]), .b(b[0]), .ci(ci), .s(s[0]));
	fa_v2 cla_fa1 (.a(a[1]), .b(b[1]), .ci(c[0]), .s(s[1]));
	fa_v2 cla_fa2 (.a(a[2]), .b(b[2]), .ci(c[1]), .s(s[2]));
	fa_v2 cla_fa3 (.a(a[3]), .b(b[3]), .ci(c[2]), .s(s[3]));
	
	clb4 clb40(.a(a), .b(b), .ci(ci), .c1(c[0]), .c2(c[1]), .c3(c[2]), .co(co));
	
endmodule
